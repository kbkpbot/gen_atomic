module main

import os
import strings
import arrays.diff
import time

// Supported CPU architectures
const archs = ['i386', 'x86_64', 'arm', 'aarch64', 'riscv']
// Atomic functions requiring size suffix (1/2/4/8 bytes)
const funcs_4 = [
	'__atomic_load',
	'__atomic_store',
	'__atomic_compare_exchange',
	'__atomic_exchange',
	'__atomic_fetch_add',
	'__atomic_add_fetch',
	'__atomic_fetch_sub',
	'__atomic_sub_fetch',
	'__atomic_fetch_and',
	'__atomic_and_fetch',
	'__atomic_fetch_or',
	'__atomic_or_fetch',
	'__atomic_fetch_nand',
	'__atomic_nand_fetch',
	'__atomic_fetch_xor',
	'__atomic_xor_fetch',
	'__atomic_test_and_set',
]

// Atomic functions not requiring size suffix
const funcs_1 = [
	'atomic_thread_fence',
	'atomic_signal_fence',
	'atomic_flag_test_and_set',
	'atomic_flag_test_and_set_explicit',
	'atomic_flag_clear',
	'atomic_flag_clear_explicit',
]

// gen_objdump_file generates disassembly output for a specific function
fn gen_objdump_file(a string, f string, need_fix bool, no_addresses bool, fix_label bool) []string {
	// Format function name for search if needed
	ff := if need_fix { 'libat_' + f.all_after('__atomic_') } else { f }

	// Execute objdump to disassemble the function
	// Note: you need an objdump which supports *ALL* archs
	mut cmd := '/usr/bin/objdump -d --disassemble=${ff} ${a}'
	if no_addresses {
		cmd = '/usr/bin/objdump -d --disassemble=${ff} --no-addresses ${a}'
	}
	result := os.execute(cmd)

	mut output := []string{}
	for line in result.output.split_into_lines() {
		// Filter out irrelevant lines
		if line.contains('.o:') || line.contains('.o：') || line.contains('libatomic.a')
			|| line.contains('Disassembly') || line.contains('>:') || line.len == 0 {
			continue
		}
		// Apply name substitution if needed
		if need_fix {
			output << line.replace('libat_', '__atomic_').expand_tabs(4).all_before(';')
		} else {
			output << line.expand_tabs(4).all_before(';')
		}
	}
	if fix_label {
		return fix_objdump_asm(output, f)
	}
	return output
}

// fix_objdump_asm fixes label formats in objdump output
fn fix_objdump_asm(src []string, f string) []string {
	mut result1 := []string{}
	mut result2 := []string{}
	mut labels := map[string]bool{} // Track found labels

	// Process each line of disassembly
	for s in src {
		if s.contains('#') {
			result1 << s
		} else if pos1 := s.index(' <') {
			// Handle jump target formatting:
			// Original: "1d <__atomic_fetch_add_8+0x1d>"
			// Convert to: ".L___atomic_fetch_add_8_1d"
			// bne t3,a7,44 <.L1^B2>
			mut pos2 := 0
			for i := pos1 - 1; i > 0; i-- {
				if s[i] in [`0`, `1`, `2`, `3`, `4`, `5`, `6`, `7`, `8`, `9`, `a`, `b`, `c`, `d`,
					`e`, `f`] {
					continue
				}
				pos2 = i + 1
				break
			}
			mut addr := s[pos2..pos1].trim_space()
			if addr.len == 1 {
				addr = '0' + addr
			} else if addr.len > 2 {
				panic('error! addr len > 2 : ${f} ${s} addr=${addr}')
			}
			result1 << s[..pos2] + ' .L_${f}_${addr}'
			labels[addr] = true // Mark as found label
		} else {
			result1 << s
		}
	}

	// Process and insert label definitions
	mut all_labels := labels.keys()
	all_labels.sort() // Sort labels for consistent ordering
	mut l := ''
	mut ss := ''
	for s in result1 {
		mut addr := s.all_before(':').trim_space()
		// Insert label definition if it matches
		if addr.len == 1 {
			addr = '0' + addr
		}
		if all_labels.len > 0 {
			l = all_labels[0]
			if l == addr {
				ss = '.L_${f}_${l}:'
				result2 << ss
				all_labels = all_labels[1..].clone() // Move to next label
			}
		}
		result2 << s
	}
	if all_labels.len > 0 {
		println('Error! lables not found for ${f}: ${all_labels}')
	}
	return result2
}

// output_global_header outputs global file header with metadata
fn output_global_header(mut sb strings.Builder) {
	sb.writeln('/* ---------------------------------------------- */')
	sb.writeln('/* This file is extracted from `gcc` v15.1.0 `libatomic.a`. */')
	sb.writeln('/* This file is generated by https://github.com/kbkpbot/gen_atomic.git */')
	now := time.now().format()
	sb.writeln('/* This file is generated at ${now}. */')
	sb.write_string('/* This file implements for ')
	sb.write_string(archs.join('/'))
	sb.writeln(':')

	// List all implemented functions
	for f in funcs_4 {
		sb.writeln(' * ${f}_[1,2,4,8]')
	}
	for f in funcs_1 {
		sb.writeln(' * ${f}')
	}
	sb.writeln(' */')

	// Handle leading underscore for symbols
	sb.writeln('#ifdef __leading_underscore')
	sb.writeln('# define _(s) _##s')
	sb.writeln('#else')
	sb.writeln('# define _(s) s')
	sb.writeln('#endif\n')
}

// output_f_header outputs function header (symbol definition)
fn output_f_header(mut sb strings.Builder, f string) {
	sb.writeln('        .global _(${f})')
	sb.writeln('        .type   _(${f}), %function')
	sb.writeln('_(${f}):')
}

// output_f_body_machine_code outputs function body as machine code instructions
fn output_f_body_machine_code(mut sb strings.Builder, f string, all []string) {
	mut c := []string{}
	for line in all {
		if line.starts_with('.L') {
			continue
		}
		ff := line.trim_space().fields()
		if ff.len > 2 {
			s := ff[1]
			if s.len == 8 {
				c << '        .int 0x' + ff[1]
			} else if s.len == 4 {
				c << '        .short 0x' + ff[1]
			} else {
				println('error! machine code line not correct: ${line}')
			}
		}
	}
	x := c.join_lines()
	sb.writeln(x)
}

// output_f_body output function body as assembly instructions
fn output_f_body(mut sb strings.Builder, f string, all []string, pos int) {
	mut c := []string{}
	for line in all {
		if line.starts_with('.L') {
			c << line
		} else {
			inst := line[pos..].trim_space()
			c << '        ' + inst
		}
	}

	x := c.join_lines()
	sb.writeln(x)
}

// output_f_footer outputs function footer (size calculation)
fn output_f_footer(mut sb strings.Builder, f string) {
	sb.writeln('	.size   _(${f}), .-_(${f})\n')
}

// output_arch_header outputs architecture-specific section header
fn output_arch_header(mut sb strings.Builder, arch string) {
	sb.writeln('\n/* ---------------------------------------------- */')
	match arch {
		'i386' {
			sb.writeln('#if defined __i386__')
		}
		'x86_64' {
			sb.writeln('#if defined __x86_64__')
		}
		'arm' {
			sb.writeln('#if defined __arm__')
		}
		'aarch64' {
			sb.writeln('#if defined __aarch64__')
		}
		'riscv' {
			sb.writeln('#if defined __riscv')
		}
		else {}
	}
	sb.writeln('        .text')
	sb.writeln('        .align  2')
	if arch == 'arm' {
		sb.writeln('        .thumb')
		sb.writeln('        .syntax unified')
	}
	sb.writeln('')
}

// output_arch_footer outputs architecture-specific section footer
fn output_arch_footer(mut sb strings.Builder, arch string) {
	match arch {
		'i386' {
			sb.writeln('#endif //__i386__')
		}
		'x86_64' {
			sb.writeln('#endif //__x86_64__')
		}
		'arm' {
			sb.writeln('#endif //__arm__')
		}
		'aarch64' {
			sb.writeln('#endif //__aarch64__')
		}
		'riscv' {
			sb.writeln('#endif //__riscv')
		}
		else {}
	}
}

// process_arch generates assembly for all functions in a specific architecture
fn process_arch(mut sb strings.Builder, arch string) ! {
	output_arch_header(mut sb, arch)

	// Architecture-specific library file
	lib_file := './libatomic.a.' + arch
	println('processing ${lib_file}...')
	mut all := []string{}
	mut need_fix := false
	// Determine disassembly format for this arch
	pos := match arch {
		'i386', 'x86_64' {
			27
		} // x86 disassembly position
		'arm', 'aarch64' {
			20
		} // ARM disassembly position
		'riscv' {
			28
		} // RISC-V disassembly position
		else {
			0
		}
	}

	mut all_funcs := []string{}
	for f in funcs_4 {
		for i in [1, 2, 4, 8] {
			all_funcs << f + '_${i}'
		}
	}
	for f in funcs_1 {
		all_funcs << f
	}

	for f in all_funcs {
		output_f_header(mut sb, f)
		need_fix = arch in ['aarch64', 'arm'] && f.starts_with('__atomic_')
		all = gen_objdump_file(lib_file, f, need_fix, false, true)
		if arch in ['riscv', 'aarch64', 'arm'] {
			sb.writeln('#ifdef __TINYC__')
			output_f_body_machine_code(mut sb, f, all)
			sb.writeln('#else')
		}
		output_f_body(mut sb, f, all, pos)
		output_f_footer(mut sb, f)
		if arch in ['riscv', 'aarch64', 'arm'] {
			sb.writeln('#endif')
		}
	}

	output_arch_footer(mut sb, arch)
}

// verify verifies generated `atomic.S` by compiling it to `atomic.o` and then verifying it with `objdump`
fn verify() {
	mut need_fix := false
	for arch in archs {
		println('verifying ${arch}')
		// Step 1: Compile atomic.S into object file
		mut cmd := ''
		lib_file := './libatomic.a.' + arch
		match arch {
			'i386' {
				cmd = '/usr/bin/i686-linux-gnu-gcc'
			}
			'x86_64' {
				cmd = '/usr/bin/gcc'
			}
			'arm' {
				cmd = '/home/mars/gcc/arm-gnu-toolchain-14.2.rel1-aarch64-arm-none-linux-gnueabihf/bin/arm-none-linux-gnueabihf-gcc'
			}
			'aarch64' {
				cmd = '/usr/bin/gcc'
			}
			'riscv' {
				cmd = '/usr/bin/gcc'
			}
			else {
				panic('unknown arch ${arch}')
			}
		}
		result := os.execute('${cmd} -c atomic.S')
		dump(cmd)
		assert result.exit_code == 0

		// Step 2: Disassemble the file using objdump
		mut all_funcs := []string{}
		for f in funcs_4 {
			for i in [1, 2, 4, 8] {
				all_funcs << f + '_${i}'
			}
		}
		for f in funcs_1 {
			all_funcs << f
		}

		for f in all_funcs {
			need_fix = arch in ['aarch64', 'arm'] && f.starts_with('__atomic_')
			orig_all := gen_objdump_file(lib_file, f, need_fix, true, false)
			new_all := gen_objdump_file('./atomic.o', f, false, true, false)
			mut df := diff.diff[string](orig_all, new_all)
			str := df.generate_patch()
			if str != '' {
				println('${arch}, ${f} :')
				println(str)
			}
		}
	}
}

fn main() {
	println('==== A libatomic.a ==> atomic.S converter for TinyCC ====')
	println('NOTE: you need an `objdump` which supports *ALL* archs')
	mut file_not_exist := false
	for arch in archs {
		f := './libatomic.a.${arch}'
		if !os.exists(f) {
			println('you need a file here: ${f}')
			file_not_exist = true
		}
	}
	if file_not_exist {
		return
	}
	mut sb := strings.new_builder(8192)

	output_global_header(mut sb)

	for arch in archs {
		process_arch(mut sb, arch)!
	}
	println('writing out atomic.S')
	os.write_file('atomic.S', sb.str())!
	// verify()
}
